** Profile: "SCHEMATIC1-sim2"  [ C:\Users\Cthulhu\Downloads\IoT_project-master\OrCAD\Amplificador_PTC\Amplificador_ptc-PSpiceFiles\SCHEMATIC1\sim2.sim ] 

** Creating circuit file "sim2.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Cthulhu\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
